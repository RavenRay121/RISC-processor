module tem(
    input a,
    output b
);
assign b = a;
endmodule